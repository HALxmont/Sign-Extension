--------------------------------------------------------------------------------
-- Company: UBB
-- Engineer: Mauricio Montanares
--
-- Create Date:   22:16:27 10/28/2018
-- Design Name:   
-- Module Name:   /home/xmont/Proyectos Git/sign extension vhdl/Sign_extension/B_signex.vhd
-- Project Name:  Sign_extension
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: sign_extension
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 

 
ENTITY B_signex IS
END B_signex;
 
ARCHITECTURE behavior OF B_signex IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT sign_extension
    PORT(
         u : IN  std_logic_vector(15 downto 0);
         y : OUT  std_logic_vector(31 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal u : std_logic_vector(15 downto 0) := (others => '0');

 	--Outputs
   signal y : std_logic_vector(31 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
   --constant <clock>_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: sign_extension PORT MAP (
          u => u,
          y => y
        );

   -- Clock process definitions
--   <clock>_process :process
--		begin
--		<clock> <= '0';
--		wait for <clock>_period/2;
--		<clock> <= '1';
--		wait for <clock>_period/2;
--   end process;
 
--		Stimulus Process
	
-- The code of below its here only for see something in simulation	
		stim_proc: process
		begin
		 
		wait for 100 ns;
		u <= x"0123";
		wait for 100 ns;
		u <= x"8123";
		wait for 100 ns;
		u <= x"F123";
		
		wait;
		end process;
END;
